library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

architecture TestBehavior of Test is
begin
  b <= a;
end architecture TestBehavior;
