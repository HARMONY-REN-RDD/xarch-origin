library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Test is
  port (
    a : in std_logic;
    b : out std_logic
  );
end entity Test;
